SAR Logic Part

.lib "./sky130.lib.spice" tt


.ic V(A)=0 V(B)=0 V(C)=0 V(D)=0 V(E)=0 V(F)=0 V(G)=0 V(H)=0 V(I)=0 V(D0_)=0 V(D1_)=0 V(D2_)=0 V(D3_)=0 V(D4_)=0 V(D5_)=0 V(D6_)=0 V(D7_)=0 V(D8_)=0 V(D9_)=0 V(dac_out)=0 V(inm)=0 V(inp)=0 V(comp__out)=0 V(V_SAM)=0 V(VIN)=0

XClk_div q0b q0 q1b q1 q2b q2 q3b q3 1 0 CLK clkdiv
Xn_o 1 0 q2 q2p q2n non_overlap
Xand 0 1 q2p q3 clk_sam1  AND_2
Xsam 1 0 VIN V_SAM clk_sam1 s_h
Xdac10 1 0 vref d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 d0_ d1_ d2_ d3_ d4_ d5_ d6_ d7_ d8_ d9_ A B C D E F G H I dac_out dac10
XSAR 1 0 CLK SOC EOC comp__out d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 SAR
Xcomp inp inm clk_preamp clk_latch om2 comp_out op1 om1 1 0 Comparator
Xinv 1 0  clk_preamp clk_latch inv
*Clock Divider
.subckt clkdiv q0b q0 q1b q1 q2b q2 q3b q3  VDD 0 CLK
XU1 0 VDD q0b 0 0 q0 q0b CLK DFFSR
XU2 0 VDD q1b 0 0 q1 q1b q0 DFFSR
XU3 0 VDD q2b 0 0 q2 q2b q1 DFFSR
XU4 0 VDD q3b 0 0 q3 q3b q2 DFFSR
.ends
*Non-Overlapping Clock Generator
.subckt non_overlap 1 0 clk1 phi1 phi2
X1 1 0 clk1 clk2 inv
X2 1 0 clk1 no2 no1 nand
X3 1 0 clk2 no1 no2 nand
X4 1 0 no1 phi1 inv
X5 1 0 no2 phi2 inv
.ends non_overlap
*Inverter
.subckt inv 1 0 in out
XM10 out in 1 1 sky130_fd_pr__pfet_01v8 W= 4 L=0.150
XM20 out in 0 0 sky130_fd_pr__nfet_01v8 W= 2.4 L=0.150
.ends inv
*NAND
.subckt nand 1 0 A B out
XM00 out A 1 1 sky130_fd_pr__pfet_01v8 W= 2 L=0.150
XM01 out B 1 1 sky130_fd_pr__pfet_01v8 W= 2 L=0.150
XM10 out A x 0 sky130_fd_pr__nfet_01v8 W= 2.2 L=0.150
XM11 x B 0 0 sky130_fd_pr__nfet_01v8 W= 2.2 L=0.150
.ends nand
*AND
.subckt AND_2 0 1 IN1 IN2  OUT1
XM1 OUT IN1 1 1 sky130_fd_pr__pfet_01v8 W= 2 L=0.150
XM2 OUT IN2 1 1 sky130_fd_pr__pfet_01v8 W= 2 L=0.150
XM4 OUT IN1 P 0 sky130_fd_pr__nfet_01v8 W= 2.2 L=0.150
XM6 P IN2 0 0 sky130_fd_pr__nfet_01v8 W=2.2 L=0.150
XM22 OUT1 OUT 1 1 sky130_fd_pr__pfet_01v8 W= 1.6 L=0.150
XM33 OUT1 OUT 0 0 sky130_fd_pr__nfet_01v8 W= 0.8 L=0.150
.ends AND_2

*Sample & Hold
.subckt s_h 1 0 VIN V_SAM CLK_A 
XM1 1 3 2 0 sky130_fd_pr__nfet_01v8 l=0.150 w=1
XC1 2 CLK_B sky130_fd_pr__cap_mim_m3_1 W=13.8 L=13.8 m=1
XM2 1 2 3 0 sky130_fd_pr__nfet_01v8 l=0.150 w=1
XC2 3 4 sky130_fd_pr__cap_mim_m3_1 W=13.u L=13.8 m=1
XMCA 4 CLK_B 1 1 sky130_fd_pr__pfet_01v8 l=0.150 w=0.650
XMCB 4 CLK_B 0 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.400
XM3 1 2 5 0 sky130_fd_pr__nfet_01v8 l=0.150 w=1
XC3 5 6 sky130_fd_pr__cap_mim_m3_1 W=13.8 L=13.8 m=2
XM12 6 CLK_B 0 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.800
XMCC CLK_B CLK_A 1 1 sky130_fd_pr__pfet_01v8 l=0.150 w=0.650
XMCD CLK_B CLK_A 0 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.400
XM4 7 CLK_A 1 1 sky130_fd_pr__pfet_01v8 l=0.150 w=0.800
XM5 7 CLK_A 6 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.450
XM8 8 7 5 5 sky130_fd_pr__pfet_01v8 l=0.200 w=0.420
XM7 8 1 9 0 sky130_fd_pr__nfet_01v8 l=0.200 w= 0.420
XM10 9 CLK_B 0 0 sky130_fd_pr__nfet_01v8 l=0.200 w=0.420
XM13 7 8 6 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.500
XM9 6 8 VIN 0 sky130_fd_pr__nfet_01v8 l=0.200 w=0.400
XM11 VIN 8 V_SAM 0 sky130_fd_pr__nfet_01v8 l=0.150 w=0.450
XCsam V_SAM 0 sky130_fd_pr__cap_mim_m3_1 W=13.8 L=13.8 m=8
.ends
Bvsam inp 0 V=V(V_SAM)
Bdac inm 0 V=V(dac_out)
Bc comp__out 0 V= V(V_SAM) > V(dac_out) && V(V_SAM)> 0.75m  && V(dac_out)>0.75m  && abs(V(V_SAM)-V(dac_out)) > 0.75m ? 1.8 : 0
.subckt buf_dac 1 0 dx dxx
XM1 dx11 dx 1 1 sky130_fd_pr__pfet_01v8 l=0.2 w=1.6
XM2 dx11 dx 0 0 sky130_fd_pr__nfet_01v8 l=0.2 w=0.8
XM3 dxx1 dx11 1 1 sky130_fd_pr__pfet_01v8 l=0.2 w=3.2
XM4 dxx1 dx11 0 0 sky130_fd_pr__nfet_01v8 l=0.2 w=1.6
XM5 dx2 dxx1 1 1 sky130_fd_pr__pfet_01v8 l=0.2 w=5.6
XM6 dx2 dxx1 0 0 sky130_fd_pr__nfet_01v8 l=0.2 w=3
XM7 dxx dx2 1 1 sky130_fd_pr__pfet_01v8 l=0.2 w=6
XM8 dxx dx2 0 0 sky130_fd_pr__nfet_01v8 l=0.2 w=3
.ends buf_dac
*DAC Switches
.SUBCKT switch data node vref 1 0
XM1 node data_bar vref 1 sky130_fd_pr__pfet_01v8 L=0.3 W=16
XM2 node data_bar 0 0 sky130_fd_pr__nfet_01v8 L=0.3 W=16
XM3 data_bar data 1 1 sky130_fd_pr__pfet_01v8 L=0.2 W=6
XM4 data_bar data 0 0 sky130_fd_pr__nfet_01v8 L=0.2 W=3
.ENDS switch
*DAC Sub-block
.subckt dac10 1 0 vref d0 d1 d2 d3 d4 d5 d6 d7 d8 d9 d0_ d1_ d2_ d3_ d4_ d5_ d6_ d7_ d8_ d9_ A B C D E F G H I out 
XC1 A 0 sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC2 A D0_ sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC3 A B  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC4 B D1_  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC5 B C  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC6 C D2_  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC7 C D  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC8 D D3_ sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC9 D E  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC10 E D4_ sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC11 E F sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC12 F D5_  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC13 F G  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC14 G D6_  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC15 G H  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC16 H D7_ sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC17 H I sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC18 I D8_ sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
XC19 I out sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=2
XC20 out D9_  sky130_fd_pr__cap_mim_m3_1 W=2.8 L=2.8 m=1
X1 D00 D0_ vref  1 0 switch
X2 D01 D1_ vref  1 0 switch
X3 D02 D2_ vref  1 0 switch
X4 D03 D3_ vref  1 0 switch
X5 D04 D4_ vref  1 0 switch
X6 D05 D5_ vref  1 0 switch
X7 D06 D6_ vref 1 0 switch
X8 D07 D7_ vref  1 0 switch
X9 D08 D8_ vref  1 0 switch
X10 D09 D9_ vref  1 0 switch
XB0 1 0 d0 d00 buf_dac
XB1 1 0 d1 d01 buf_dac
XB2 1 0 d2 d02 buf_dac
XB3 1 0 d3 d03 buf_dac
XB4 1 0 d4 d04 buf_dac
XB5 1 0 d5 d05 buf_dac
XB6 1 0 d6 d06 buf_dac
XB7 1 0 d7 d07 buf_dac
XB8 1 0 d8 d08 buf_dac
XB9 1 0 d9 d09 buf_dac
.ends dac10
.subckt Comparator inp inm clk_preamp clk_latch op2 om2 op1 om1 vdd gnd
Xpreamp inp inm clk_preamp op1 om1 vdd 0 preamp
Xstrong_arm_latch om1 op1  clk_latch op2 om2 vdd 0 strong_arm_latch
.ends Comparator
.subckt preamp inp inn clk_pre opp1 opn1 1 0
XM1 2 clk_pre 1 1 sky130_fd_pr__pfet_01v8 L=2 W=1
XM2 opp1 inn 2 1 sky130_fd_pr__pfet_01v8 L=0.5 W=2
XM3 opn1 inp 2 1 sky130_fd_pr__pfet_01v8 L=0.5 W=2
XM4 opp1 clk_pre opn1 1 sky130_fd_pr__pfet_01v8 L=0.5 W=1
XM5 opp1 opp1 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=0.5
XM6 opp1 opn1 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=0.5
XM7 opn1 opp1 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=0.5
XM8 opn1 opn1 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=0.5
.ends preamp
.subckt strong_arm_latch opp1 opn1 clk_latch opp2 opn2 1 0
XM1 2 clk_latch 1 1 sky130_fd_pr__pfet_01v8 L=1 W=24
XM2 3 opn1 2 1 sky130_fd_pr__pfet_01v8 L=0.35 W=12
XM3 4 opp1 2 1 sky130_fd_pr__pfet_01v8 L=0.35 W=12
XM4 opp2 opn2 3 1 sky130_fd_pr__pfet_01v8 L=0.35 W=6
XM5 opn2 opp2 4 1 sky130_fd_pr__pfet_01v8 L=0.35 W=6
XM6 opp2 opn2 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=3
XM7 opp2 clk_latch 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=3
XM8 opn2 opp2 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=3
XM9 opn2 clk_latch 0 0 sky130_fd_pr__nfet_01v8 L=0.5 W=3
.ends strong_arm_latch 
.subckt SAR VDD 0 CLK SOC EOC COMP D0 D1 D2 D3 D4 D5 D6 D7 D8 D9
XU1 0 VDD 0 SOC 0 q1 q1b CLK DFFSR
XU2 0 VDD q1 0 SOC q2 q2b CLK DFFSR
XU3 0 VDD q2 0 SOC q3 q3b CLK DFFSR
XU4 0 VDD q3 0 SOC q4 q4b CLK DFFSR
XU5 0 VDD q4 0 SOC q5 q5b CLK DFFSR
XU6 0 VDD q5 0 SOC q6 q6b CLK DFFSR
XU7 0 VDD q6 0 SOC q7 q7b CLK DFFSR
XU8 0 VDD q7 0 SOC q8 q8b CLK DFFSR
XU9 0 VDD q8 0 SOC q9 q9b CLK DFFSR
XU10 0 VDD q9 0 SOC q10 q10b CLK DFFSR
XU11 0 VDD q10 0 SOC EOC q11b CLK DFFSR
XU12 0 VDD 0 EOC SOC q12 q12b 0 DFFSR
XU13 0 VDD COMP q10 SOC d0 d0b q12 DFFSR
XU14 0 VDD COMP q9 SOC d1 d1b d0 DFFSR
XU15 0 VDD COMP q8 SOC d2 d2b d1 DFFSR
XU16 0 VDD COMP q7 SOC d3 d3b d2 DFFSR
XU17 0 VDD COMP q6 SOC d4 d4b d3 DFFSR
XU18 0 VDD COMP q5 SOC d5 d5b d4 DFFSR
XU19 0 VDD COMP q4 SOC d6 d6b d5 DFFSR
XU20 0 VDD COMP q3 SOC d7 d7b d6 DFFSR
XU21 0 VDD COMP q2 SOC d8 d8b d7 DFFSR
XU22 0 VDD COMP q1 SOC d9 d9b d8 DFFSR
.ends SAR
.subckt DFFSR 0 1 D S R Q Q_bar CLK
XM1 2 D 1 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM2 3 CLK 2 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM3 3 D 0 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM4 4 CLK 1 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM5 4 3 5 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM6 5 CLK 0 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM7 6 4 1 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM8 6 CLK 7 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM9 7 4 0 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM10 6 R_bar 1 1 sky130_fd_pr__pfet_01v8 W= 1.6 L=0.150
XM11 6 S 0 0 sky130_fd_pr__nfet_01v8 W=0.800 L=0.150
XM12 R_bar R 1 1 sky130_fd_pr__pfet_01v8 W= 1.6 L=0.150
XM13 R_bar R 0 0 sky130_fd_pr__nfet_01v8 W= 0.800 L=0.150
XM14 Q 6 1 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM15 Q 6 0 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
XM16 Q_bar Q 1 1 sky130_fd_pr__pfet_01v8 W= 0.600 L=0.150
XM17 Q_bar Q 0 0 sky130_fd_pr__nfet_01v8 W= 0.400 L=0.150
.ends DFFSR
*______________________________________________________________

BV9 b9 0 V= V(d9)>1.5 ? 1 : 0
BV8 b8 0 V= V(d8)>1.5 ? 1 : 0
BV7 b7 0 V= V(d7)>1.5 ? 1 : 0
BV6 b6 0 V= V(d6)>1.5 ? 1 : 0
BV5 b5 0 V= V(d5)>1.5 ? 1 : 0
BV4 b4 0 V= V(d4)>1.5 ? 1 : 0
BV3 b3 0 V= V(d3)>1.5 ? 1 : 0
BV2 b2 0 V= V(d2)>1.5 ? 1 : 0
BV1 b1 0 V= V(d1)>1.5 ? 1 : 0
BV0 b0 0 V= V(d0)>1.5 ? 1 : 0
BVc code 0 V= V(b9)*512 + V(b8)*256 + V(b7)*128 + V(b6)*64 + V(b5)*32 + V(b4)*16 + V(b3)*8 + V(b2)*4 + V(b1)*2 + V(b0)*1
BVa analog 0 V= 0.001757*V(code)
*______________________________________________________________
****************************************************************************************
*V9 D9 0 PULSE(1.8V 0 1p 1p 1p 12800n 25600n)
*V8 D8 0 PULSE(1.8V 0 1p 1p 1p 6400n 12800n)
*V7 D7 0 PULSE(1.8V 0 1p 1p 1p 3200n 6400n)
*V6 D6 0 PULSE(1.8V 0 1p 1p 1p 1600n 3200n)
*V5 D5 0 PULSE(1.8V 0 1p 1p 1p 800n 1600n)
*V4 D4 0 PULSE(1.8V 0 1p 1p 1p 400n 800n)
*V3 D3 0 PULSE(1.8V 0 1p 1p 1p 200n 400n)
*V2 D2 0 PULSE(1.8V 0 1p 1p 1p 100n 200n)
*V1 D1 0 PULSE(1.8V 0 1p 1p 1p 50n 100n)
*V0 D0 0 PULSE(1.8V 0 1p 1p 1p 25n 50n)
Vsoc SOC 0 PULSE(0 1.8 200n 1n 1n 0.028u 0.8u)
Vclk CLK 0 PULSE(0 1.8 1p 1p 1p 0.025u 0.05u)
Vclk1 clk_preamp  0 PULSE(1.8 0 0.0125u 1p 1p 0.025u 0.05u )

*__________________________INPUT HERE______________________________________



BVI VIN 0 V= 393.75*time + 1.564614125


Vdd 1 0 dc 1.8
Vd_vref vref 0 1.8

.control
*************************************************************************
set num_threads=8
*************************************************************************
run

tran 0.001u 662u 0us
let ideal = V(V_SAM)/0.001757
let lin-tstart =1.57us
let lin-tstop=662us
let lin-tstep=0.8us
linearize V_SAM code ideal


print time V_SAM code > ./DATA/final8.csv 


.endc
.end


